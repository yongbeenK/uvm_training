// apb_top
module top

// dut
// env
// clock
// interface
// run_test();

endmodule
