// APB test

class apb_test extends uvm_test

endclass
