// top

module top

// clock
// interface
//  run_test();

endmodule
