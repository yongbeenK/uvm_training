// apb_incr_top.sv
module incr_top

// for changeable thing
// interface

endmodule
