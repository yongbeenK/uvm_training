// top

module top



endmoudle
