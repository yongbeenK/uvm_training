// apb_dut - buffer or inverter
module dut

endmodule
