
interface buffer_intf 
  logic a;
  logic b;
  logic en;

endinterface
