// apb_top
module top

// dut
  apb_dut apb_test_dut_0();
// env
// clock
// interface
// run_test();

endmodule
